`define GLOBAL_BUSADDRWID 32
`define GLOBAL_BUSDATAWID 64
`define GPU_DDATA_WIDTH 32
`define GPU_DADDR_WIDTH 32
`define GPU_IADDR_WIDTH 32
`define GPU_VDATA_WIDTH `GPU_LANE_WIDTH*GPU_LANE_NUM
`define GPU_LANE_WIDTH 16
`define GPU_LANE_NUM 8

