module backend_top
(
);





endmodule
