module GPR
(
    input [4:0]rs1,
    input [4:0]rs2,
    output [31:0]rs1o,
    output [31:0]rs2o,
    input [31:0]rdi,
    input [4:0]rd,
    input rdw,
    input clk
);
reg [31:0]regs[31:1];
assign rs1o=(rs1==0)?32'b0:regs[rs1];
assign rs2o=(rs2==0)?32'b0:regs[rs2];
always @(posedge clk)
begin
    if(rdw&rd!=0)
        regs[rd]<=rdi;
end

endmodule