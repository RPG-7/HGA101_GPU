`define GLOBAL_BUSADDRWID 32
`define GLOBAL_BUSDATAWID 32
`define FCU_DDATA_WIDTH 32
`define FCU_IADDR_WIDTH 32



