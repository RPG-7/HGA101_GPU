`define GLOBAL_BUSADDRWID 64
`define GLOBAL_BUSDATAWID 64
`define GPU_CACHE_DATAWID 64
`define GPU_DDATA_WIDTH 64
`define GPU_DADDR_WIDTH 64
`define GPU_IADDR_WIDTH 64

`define GPU_LANE_WIDTH 16
`define GPU_LANE_NUM 8

`define GPU_VDATA_WIDTH `GPU_LANE_WIDTH*`GPU_LANE_NUM
`define DUMP_VCD