module fpu32
(
    
);




endmodule
