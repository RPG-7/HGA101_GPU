module CORDIC16
();




endmodule
